module sdram_write(

);

endmodule
