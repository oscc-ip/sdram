module clk();

endmodule
