`timescale 1ns / 1ns;

module tb_clk();

endmodule
