`timescale  1ns / 1ns;

module tb_sdram_fifo();

endmodule
