module axi4(

);

endmodule
